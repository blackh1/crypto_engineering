`timescale 1ns/1ps

module cipher(clk,msg,pubk,prik,out,ans);


always @(posedge clk)
begin

end